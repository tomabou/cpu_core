module hazard_detect