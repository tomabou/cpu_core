module ip_test();

endmodule
