module int_to_float();

endmodule
