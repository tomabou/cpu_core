module nibu (clk);
    input clk;

endmodule