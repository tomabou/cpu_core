module akari(clk,rxd,seg1,seg2,seg3,seg4,seg5,seg6,txd);
    input clk;
    input rxd;
    output [6:0] seg1;
    output [6:0] seg2;
    output [6:0] seg3;
    output [6:0] seg4;
    output [6:0] seg5;
    output [6:0] seg6;
    output txd;
    wire slow_clk;

endmodule

