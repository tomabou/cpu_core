module float_to_int(
    x,
    is_cvt,
    y);
    input [31:0] x;
    input is_cvt;
    output [31:0] y;

    assign y = x;

endmodule
