module fpu_control();

endmodule
