module forward_ctl ()