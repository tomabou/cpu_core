module uart_input(clk,input);
