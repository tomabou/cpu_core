module akari();

endmodule

