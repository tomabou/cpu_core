module float_to_int();

endmodule
